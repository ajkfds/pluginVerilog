`timescale 1n/1p

module DIMENSIONS;

wire [7:0] a [0:10];
wire [7:0] b;


assign	a[1][0] = b[1];
assign	a[1][0] = b[1];
	assign	a[1][0] = b[1];
	assign	a[1][0] = b[1];



endmodule