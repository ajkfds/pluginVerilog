module MOD3(
input	CLK_I,
input	RST_X
);



endmodule
endmo