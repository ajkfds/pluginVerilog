module REAL_CONSTANTS;


// Examples:


real r0 = 1.2;

real r1 = 0.1;
real r2 = 394.26331;
real r3 = 1.2E12; // (the exponent symbol can be e or E)
real r4 = 1.30e-2;
real r5 = 0.1e-0;
real r6 = 23E10;
real r7 = 29E-2;
real r8 = 236.123_763_e-12;//  (underscores are ignored)
//The following are invalid forms of real numbers because they do not have at least one digit on each side of the decimal point:
real r9 = .12;
real r10 9. 
 4.E3 
 .2e-7

endmodule
