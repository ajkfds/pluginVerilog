
module MOD(
output [7:0]	DATA_O,
input	CLK_I,
inout aaa,
input	RST_X
);

assign DATA_O = 8'h01;
reg [7:0] regMod;


endmodule


endmodule