
module TEST_TOP3;


TOP #(
	.WIDTH	(  )
)  TOP_0 (
	.DATA_I	(  ),
	.DATA_O	(  ),
	.CLK_I	(  ),
	.RST_X	(  )
);


endmodule


