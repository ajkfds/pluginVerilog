
localparam P_BLANK = 8'h00;
